module microcode(
    input [9:0] addr,
    output [17:0] data
);

endmodule
